module InvMixColumns(data_in, data_out);
input [127:0] data_in;
output [127:0] data_out;

GaloisMulti invmixcolumns(128'h0E090D0B0B0E090D0D0B0E09090D0B0E, data_in, data_out);

endmodule